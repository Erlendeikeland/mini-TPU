library ieee;
use ieee.std_logic_1164.all;

entity axi_tb is
end entity axi_tb;

architecture behave of axi_tb is

    

begin

    

end architecture;