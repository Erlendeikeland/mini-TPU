library ieee;
use ieee.std_logic_1164.all;

entity pe_tb is
end entity pe_tb;

architecture behave of pe_tb is

begin

    

end architecture;