library ieee;
use ieee.std_logic_1164.all;

use work.minitpu_pkg.all;

entity tpu is
    port (
        clk : in std_logic;
        reset : in std_logic

    );
end entity tpu;

architecture behave of tpu is

    

begin

    

end architecture;