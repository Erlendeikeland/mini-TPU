library ieee;
use ieee.std_logic_1164.all;

use work.minitpu_pkg.all;

entity accumulator is
    port (
        clk : in std_logic;
        
    );
end entity accumulator;

architecture behave of accumulator is

begin

    

end architecture;